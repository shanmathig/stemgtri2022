module OR2 #() (
	input wire a,
	input wire b,
	output wire o
	);

	assign o = a || b;

endmodule
