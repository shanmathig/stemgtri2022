module AND3 #() (
	input wire a,
	input wire b,
	input wire c,
	output wire o
	);

	assign o = a && b && c;

endmodule
