module INV #() (
	input wire a,
	output wire o
	);

	assign o = ~a;

endmodule
